
-- Code Store ROM

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-- USE IEEE.numeric_std.all;
use IEEE.math_real.all;
use ieee.std_logic_arith.all;
 
entity code_store_rom is
generic(
    address_length: natural := 9;
    data_length: natural := 36
);
port(
		start_signal: in std_logic;
		clock: in std_logic;
    address: in std_logic_vector((address_length - 1) downto 0);
    data_output: out std_logic_vector ((data_length - 1) downto 0)
);
end entity code_store_rom;
 
architecture a_code_store_rom of code_store_rom is
    type rom_type is array (0 to (2**(address_length) -1)) of std_logic_vector((data_length - 1) downto 0);
    
    -- set the data on each adress to some value)
    constant mem: rom_type:=
    (
			"000000001000100001000010011010000000",	-- 0 - 0
			"000000010001100100000000000001000000",	-- 1 - 1
			"000000000001001000000000000000000010",	-- 2 - 2
			"000000000000000000000000000000000000",	-- 3 - 3
			"000000000000000000000000000000000000",	-- 4 - 4
			"000000000000000000000000000000000000",	-- 5 - 5
			"000000000000000000000000000000000000",	-- 6 - 6
			"000000000000000000000000000000000000",	-- 7 - 7
			"000000000000000000000000000000000000",	-- 10 - 8
			"000000000000000000000000000000000000",	-- 11 - 9
			"000000000000000000000000000000000000",	-- 12 - 10
			"000000000000000000000000000000000000",	-- 13 - 11
			"000000000000000000000000000000000000",	-- 14 - 12
			"000000000000000000000000000000000000",	-- 15 - 13
			"000000000000000000000000000000000000",	-- 16 - 14
			"000000000000000000000000000000000000",	-- 17 - 15
			"000000000000000000000000000000000000",	-- 20 - 16
			"000000000000000000000000000000000000",	-- 21 - 17
			"000000000000000000000000000000000000",	-- 22 - 18
			"000000000000000000000000000000000000",	-- 23 - 19
			"000000000000000000000000000000000000",	-- 24 - 20
			"000000000000000000000000000000000000",	-- 25 - 21
			"000000000000000000000000000000000000",	-- 26 - 22
			"000000000000000000000000000000000000",	-- 27 - 23
			"000000000000000000000000000000000000",	-- 30 - 24
			"000000000000000000000000000000000000",	-- 31 - 25
			"000000000000000000000000000000000000",	-- 32 - 26
			"000000000000000000000000000000000000",	-- 33 - 27
			"000000000000000000000000000000000000",	-- 34 - 28
			"000000000000000000000000000000000000",	-- 35 - 29
			"000000000000000000000000000000000000",	-- 36 - 30
			"000000000000000000000000000000000000",	-- 37 - 31
			"000000000000000000000000000000000000",	-- 40 - 32
			"000000000000000000000000000000000000",	-- 41 - 33
			"000000000000000000000000000000000000",	-- 42 - 34
			"000000000000000000000000000000000000",	-- 43 - 35
			"000000000000000000000000000000000000",	-- 44 - 36
			"000000000000000000000000000000000000",	-- 45 - 37
			"000000000000000000000000000000000000",	-- 46 - 38
			"000000000000000000000000000000000000",	-- 47 - 39
			"000000000000000000000000000000000000",	-- 50 - 40
			"000000000000000000000000000000000000",	-- 51 - 41
			"000000000000000000000000000000000000",	-- 52 - 42
			"000000000000000000000000000000000000",	-- 53 - 43
			"000000000000000000000000000000000000",	-- 54 - 44
			"000000000000000000000000000000000000",	-- 55 - 45
			"000000000000000000000000000000000000",	-- 56 - 46
			"000000000000000000000000000000000000",	-- 57 - 47
			"000000000000000000000000000000000000",	-- 60 - 48
			"000000000000000000000000000000000000",	-- 61 - 49
			"000000000000000000000000000000000000",	-- 62 - 50
			"000000000000000000000000000000000000",	-- 63 - 51
			"000000000000000000000000000000000000",	-- 64 - 52
			"000000000000000000000000000000000000",	-- 65 - 53
			"000000000000000000000000000000000000",	-- 66 - 54
			"000000000000000000000000000000000000",	-- 67 - 55
			"000000000000000000000000000000000000",	-- 70 - 56
			"000000000000000000000000000000000000",	-- 71 - 57
			"000000000000000000000000000000000000",	-- 72 - 58
			"000000000000000000000000000000000000",	-- 73 - 59
			"000000000000000000000000000000000000",	-- 74 - 60
			"000000000000000000000000000000000000",	-- 75 - 61
			"000000000000000000000000000000000000",	-- 76 - 62
			"000000000000000000000000000000000000",	-- 77 - 63
			"010000000010000000010000000000000100",	-- 100 - 64
			"000000000000000000000000000000000000",	-- 101 - 65
			"000000000000000000000000000000000000",	-- 102 - 66
			"000000000000000000000000000000000000",	-- 103 - 67
			"000000000000000000000000000000000000",	-- 104 - 68
			"000000000000000000000000000000000000",	-- 105 - 69
			"000000000000000000000000000000000000",	-- 106 - 70
			"000000000000000000000000000000000000",	-- 107 - 71
			"001001001010000001000000010001000000",	-- 110 - 72
			"010000000001000000010000000000000100",	-- 111 - 73
			"000000000000000000000000000000000000",	-- 112 - 74
			"000000000000000000000000000000000000",	-- 113 - 75
			"000000000000000000000000000000000000",	-- 114 - 76
			"000000000000000000000000000000000000",	-- 115 - 77
			"000000000000000000000000000000000000",	-- 116 - 78
			"000000000000000000000000000000000000",	-- 117 - 79
			"001010001010000001000010011010000000",	-- 120 - 80
			"001010010001110000000000000001000011",	-- 121 - 81
			"001010011001000001000000010001000000",	-- 122 - 82
			"010000000001000000010000000000000100",	-- 123 - 83
			"000000000000000000000000000000000000",	-- 124 - 84
			"000000000000000000000000000000000000",	-- 125 - 85
			"000000000000000000000000000000000000",	-- 126 - 86
			"000000000000000000000000000000000000",	-- 127 - 87
			"000000000000000000000000000000000000",	-- 130 - 88
			"000000000000000000000000000000000000",	-- 131 - 89
			"000000000000000000000000000000000000",	-- 132 - 90
			"000000000000000000000000000000000000",	-- 133 - 91
			"000000000000000000000000000000000000",	-- 134 - 92
			"000000000000000000000000000000000000",	-- 135 - 93
			"000000000000000000000000000000000000",	-- 136 - 94
			"000000000000000000000000000000000000",	-- 137 - 95
			"001100001010000000000011001010000000",	-- 140 - 96
			"001100010001110001000000010001000011",	-- 141 - 97
			"001100011001000001000000010001000000",	-- 142 - 98
			"010000000001000000010000000000000100",	-- 143 - 99
			"000000000000000000000000000000000000",	-- 144 - 100
			"000000000000000000000000000000000000",	-- 145 - 101
			"000000000000000000000000000000000000",	-- 146 - 102
			"000000000000000000000000000000000000",	-- 147 - 103
			"000000000000000000000000000000000000",	-- 150 - 104
			"000000000000000000000000000000000000",	-- 151 - 105
			"000000000000000000000000000000000000",	-- 152 - 106
			"000000000000000000000000000000000000",	-- 153 - 107
			"000000000000000000000000000000000000",	-- 154 - 108
			"000000000000000000000000000000000000",	-- 155 - 109
			"000000000000000000000000000000000000",	-- 156 - 110
			"000000000000000000000000000000000000",	-- 157 - 111
			"001110001000100001000010011010000000",	-- 160 - 112
			"001110010001100100000000000001000000",	-- 161 - 113
			"001110011001000000000000000000110000",	-- 162 - 114
			"001110100010000000000010000100000000",	-- 163 - 115
			"001110110001100001000000010001000011",	-- 164 - 116
			"000000000000000000000000000000000000",	-- 165 - 117
			"001110111001000001000000010001000000",	-- 166 - 118
			"010000000001000000010000000000000100",	-- 167 - 119
			"000000000000000000000000000000000000",	-- 170 - 120
			"000000000000000000000000000000000000",	-- 171 - 121
			"000000000000000000000000000000000000",	-- 172 - 122
			"000000000000000000000000000000000000",	-- 173 - 123
			"000000000000000000000000000000000000",	-- 174 - 124
			"000000000000000000000000000000000000",	-- 175 - 125
			"000000000000000000000000000000000000",	-- 176 - 126
			"000000000000000000000000000000000000",	-- 177 - 127
			"011000000010100000100000000000110110",	-- 200 - 128
			"000000000000000000000000000000000000",	-- 201 - 129
			"000000000000000000000000000000000000",	-- 202 - 130
			"000000000000000000000000000000000000",	-- 203 - 131
			"000000000000000000000000000000000000",	-- 204 - 132
			"000000000000000000000000000000000000",	-- 205 - 133
			"000000000000000000000000000000000000",	-- 206 - 134
			"000000000000000000000000000000000000",	-- 207 - 135
			"010001001010100001000000010001000000",	-- 210 - 136
			"011000000001000000100000000000110110",	-- 211 - 137
			"000000000000000000000000000000000000",	-- 212 - 138
			"000000000000000000000000000000000000",	-- 213 - 139
			"000000000000000000000000000000000000",	-- 214 - 140
			"000000000000000000000000000000000000",	-- 215 - 141
			"000000000000000000000000000000000000",	-- 216 - 142
			"000000000000000000000000000000000000",	-- 217 - 143
			"010010001010100001000010011010000000",	-- 220 - 144
			"010010010001110100000000000001000101",	-- 221 - 145
			"010010011001000001000000010001000000",	-- 222 - 146
			"011000000001000000100000000000110110",	-- 223 - 147
			"000000000000000000000000000000000000",	-- 224 - 148
			"000000000000000000000000000000000000",	-- 225 - 149
			"000000000000000000000000000000000000",	-- 226 - 150
			"000000000000000000000000000000000000",	-- 227 - 151
			"000000000000000000000000000000000000",	-- 230 - 152
			"000000000000000000000000000000000000",	-- 231 - 153
			"000000000000000000000000000000000000",	-- 232 - 154
			"000000000000000000000000000000000000",	-- 233 - 155
			"000000000000000000000000000000000000",	-- 234 - 156
			"000000000000000000000000000000000000",	-- 235 - 157
			"000000000000000000000000000000000000",	-- 236 - 158
			"000000000000000000000000000000000000",	-- 237 - 159
			"010100001010100000000011001010000000",	-- 240 - 160
			"010100010001110101000000010001000101",	-- 241 - 161
			"010100011001000001000000010001000000",	-- 242 - 162
			"011000000001000000100000000000110110",	-- 243 - 163
			"000000000000000000000000000000000000",	-- 244 - 164
			"000000000000000000000000000000000000",	-- 245 - 165
			"000000000000000000000000000000000000",	-- 246 - 166
			"000000000000000000000000000000000000",	-- 247 - 167
			"000000000000000000000000000000000000",	-- 250 - 168
			"000000000000000000000000000000000000",	-- 251 - 169
			"000000000000000000000000000000000000",	-- 252 - 170
			"000000000000000000000000000000000000",	-- 253 - 171
			"000000000000000000000000000000000000",	-- 254 - 172
			"000000000000000000000000000000000000",	-- 255 - 173
			"000000000000000000000000000000000000",	-- 256 - 174
			"000000000000000000000000000000000000",	-- 257 - 175
			"010110001000100001000010011010000000",	-- 260 - 176
			"010110010001100100000000000001000000",	-- 261 - 177
			"010110011001000000000000000000110000",	-- 262 - 178
			"010110100010100000000010000100000000",	-- 263 - 179
			"010110110001100001000000010001000101",	-- 264 - 180
			"000000000000000000000000000000000000",	-- 265 - 181
			"010110111001000001000000010001000000",	-- 266 - 182
			"011000000001000000100000000000110110",	-- 267 - 183
			"000000000001110100000000000000000001",	-- 270 - 184
			"000000000001100010000000100001000001",	-- 271 - 185
			"000000000000000000000000000000000000",	-- 272 - 186
			"000000000000000000000000000000000000",	-- 273 - 187
			"000000000000000000000000000000000000",	-- 274 - 188
			"000000000000000000000000000000000000",	-- 275 - 189
			"000000000000000000000000000000000000",	-- 276 - 190
			"000000000000000000000000000000000000",	-- 277 - 191
			"010111000100001100000010000100000111",	-- 300 - 192
			"010111000100001100000010000000000111",	-- 301 - 193
			"010111000100001100000011000100000111",	-- 302 - 194
			"010111000100001100000011000000000111",	-- 303 - 195
			"010111000100001100000100000000000111",	-- 304 - 196
			"010111000100001100000101000000000111",	-- 305 - 197
			"010111000100001100000110000000000111",	-- 306 - 198
			"000000000100001100000011000100000001",	-- 307 - 199
			"010111000100000000000001000000000111",	-- 310 - 200
			"000000000000000000000000000000000000",	-- 311 - 201
			"000000000000000000000000000000000000",	-- 312 - 202
			"000000000000000000000000000000000000",	-- 313 - 203
			"000000000000000000000000000000000000",	-- 314 - 204
			"000000000000000000000000000000000000",	-- 315 - 205
			"000000000000000000000000000000000000",	-- 316 - 206
			"000000000000000000000000000000000000",	-- 317 - 207
			"010111000100101100000010001010000111",	-- 320 - 208
			"010111000000001100000111000000000111",	-- 321 - 209
			"010111000000001100001001000000000111",	-- 322 - 210
			"010111000000001100001010000000000111",	-- 323 - 211
			"010111000000001100001011000000000111",	-- 324 - 212
			"010111000000001100001100000000000111",	-- 325 - 213
			"010111000000001100001101000000000111",	-- 326 - 214
			"010111000000001100001110000000000111",	-- 327 - 215
			"010111000000000000001000000000000111",	-- 330 - 216
			"000000000000000000000000000000000000",	-- 331 - 217
			"000000000000000000000000000000000000",	-- 332 - 218
			"000000000000000000000000000000000000",	-- 333 - 219
			"000000000000000000000000000000000000",	-- 334 - 220
			"000000000000000000000000000000000000",	-- 335 - 221
			"000000000000000000000000000000000000",	-- 336 - 222
			"000000000000000000000000000000000000",	-- 337 - 223
			"000000000000000000000000000000000000",	-- 340 - 224
			"000000000000000000000000000000000000",	-- 341 - 225
			"000000000000000000000000000000000000",	-- 342 - 226
			"000000000000000000000000000000000000",	-- 343 - 227
			"000000000000000000000000000000000000",	-- 344 - 228
			"000000000000000000000000000000000000",	-- 345 - 229
			"000000000000000000000000000000000000",	-- 346 - 230
			"000000000000000000000000000000000000",	-- 347 - 231
			"000000000000000000000000000000000000",	-- 350 - 232
			"000000000000000000000000000000000000",	-- 351 - 233
			"000000000000000000000000000000000000",	-- 352 - 234
			"000000000000000000000000000000000000",	-- 353 - 235
			"000000000000000000000000000000000000",	-- 354 - 236
			"000000000000000000000000000000000000",	-- 355 - 237
			"000000000000000000000000000000000000",	-- 356 - 238
			"000000000000000000000000000000000000",	-- 357 - 239
			"000000000000000000000000000000000000",	-- 360 - 240
			"000000000000000000000000000000000000",	-- 361 - 241
			"000000000000000000000000000000000000",	-- 362 - 242
			"000000000000000000000000000000000000",	-- 363 - 243
			"000000000000000000000000000000000000",	-- 364 - 244
			"000000000000000000000000000000000000",	-- 365 - 245
			"000000000000000000000000000000000000",	-- 366 - 246
			"000000000000000000000000000000000000",	-- 367 - 247
			"000000000000000000000000000000000000",	-- 370 - 248
			"000000000000000000000000000000000000",	-- 371 - 249
			"000000000000000000000000000000000000",	-- 372 - 250
			"000000000000000000000000000000000000",	-- 373 - 251
			"000000000000000000000000000000000000",	-- 374 - 252
			"000000000000000000000000000000000000",	-- 375 - 253
			"000000000000000000000000000000000000",	-- 376 - 254
			"000000000000000000000000000000000000",	-- 377 - 255
			"100001000000000000000000000000001000",	-- 400 - 256
			"000000000000000000000000000000000000",	-- 401 - 257
			"000000000000000000000000000000000000",	-- 402 - 258
			"000000000000000000000000000000000000",	-- 403 - 259
			"000000000000000000000000000000000000",	-- 404 - 260
			"000000000000000000000000000000000000",	-- 405 - 261
			"000000000000000000000000000000000000",	-- 406 - 262
			"000000000000000000000000000000000000",	-- 407 - 263
			"000000000000000000000000000000000001",	-- 410 - 264
			"000000000000000000000000000000000000",	-- 411 - 265
			"000000000000000000000000000000000000",	-- 412 - 266
			"000000000000000000000000000000000000",	-- 413 - 267
			"000000000000000000000000000000000000",	-- 414 - 268
			"000000000000000000000000000000000000",	-- 415 - 269
			"000000000000000000000000000000000000",	-- 416 - 270
			"000000000000000000000000000000000000",	-- 417 - 271
			"000000000000000000000000000000000000",	-- 420 - 272
			"000000000000000000000000000000000000",	-- 421 - 273
			"000000000000000000000000000000000000",	-- 422 - 274
			"000000000000000000000000000000000000",	-- 423 - 275
			"000000000000000000000000000000000000",	-- 424 - 276
			"000000000000000000000000000000000000",	-- 425 - 277
			"000000000000000000000000000000000000",	-- 426 - 278
			"000000000000000000000000000000000000",	-- 427 - 279
			"100011001000100000000000000000110000",	-- 430 - 280
			"100011010101000000000010000100000000",	-- 431 - 281
			"000000000001100100000000000000000001",	-- 432 - 282
			"000000000000000000000000000000000000",	-- 433 - 283
			"000000000000000000000000000000000000",	-- 434 - 284
			"000000000000000000000000000000000000",	-- 435 - 285
			"000000000000000000000000000000000000",	-- 436 - 286
			"000000000000000000000000000000000000",	-- 437 - 287
			"000000000000000000000000000000000000",	-- 440 - 288
			"000000000000000000000000000000000000",	-- 441 - 289
			"000000000000000000000000000000000000",	-- 442 - 290
			"000000000000000000000000000000000000",	-- 443 - 291
			"000000000000000000000000000000000000",	-- 444 - 292
			"000000000000000000000000000000000000",	-- 445 - 293
			"000000000000000000000000000000000000",	-- 446 - 294
			"000000000000000000000000000000000000",	-- 447 - 295
			"000000000000000000000000000000000000",	-- 450 - 296
			"000000000000000000000000000000000000",	-- 451 - 297
			"000000000000000000000000000000000000",	-- 452 - 298
			"000000000000000000000000000000000000",	-- 453 - 299
			"000000000000000000000000000000000000",	-- 454 - 300
			"000000000000000000000000000000000000",	-- 455 - 301
			"000000000000000000000000000000000000",	-- 456 - 302
			"000000000000000000000000000000000000",	-- 457 - 303
			"000000000000000000000000000000000000",	-- 460 - 304
			"000000000000000000000000000000000000",	-- 461 - 305
			"000000000000000000000000000000000000",	-- 462 - 306
			"000000000000000000000000000000000000",	-- 463 - 307
			"000000000000000000000000000000000000",	-- 464 - 308
			"000000000000000000000000000000000000",	-- 465 - 309
			"000000000000000000000000000000000000",	-- 466 - 310
			"000000000000000000000000000000000000",	-- 467 - 311
			"000000000000000000000000000000000000",	-- 470 - 312
			"000000000000000000000000000000000000",	-- 471 - 313
			"000000000000000000000000000000000000",	-- 472 - 314
			"000000000000000000000000000000000000",	-- 473 - 315
			"000000000000000000000000000000000000",	-- 474 - 316
			"000000000000000000000000000000000000",	-- 475 - 317
			"000000000000000000000000000000000000",	-- 476 - 318
			"000000000000000000000000000000000000",	-- 477 - 319
			"000000000000000000000000000000001001",	-- 500 - 320
			"000000000000000000000000000000000000",	-- 501 - 321
			"000000000000000000000000000000000000",	-- 502 - 322
			"000000000000000000000000000000000000",	-- 503 - 323
			"000000000000000000000000000000000000",	-- 504 - 324
			"000000000000000000000000000000000000",	-- 505 - 325
			"000000000000000000000000000000000000",	-- 506 - 326
			"000000000000000000000000000000000000",	-- 507 - 327
			"000000000000000000000000000000000001",	-- 510 - 328
			"000000000000000000000000000000000000",	-- 511 - 329
			"000000000000000000000000000000000000",	-- 512 - 330
			"000000000000000000000000000000000000",	-- 513 - 331
			"000000000000000000000000000000000000",	-- 514 - 332
			"000000000000000000000000000000000000",	-- 515 - 333
			"000000000000000000000000000000000000",	-- 516 - 334
			"000000000000000000000000000000000000",	-- 517 - 335
			"000000000000000000000000000000000000",	-- 520 - 336
			"000000000000000000000000000000000000",	-- 521 - 337
			"000000000000000000000000000000000000",	-- 522 - 338
			"000000000000000000000000000000000000",	-- 523 - 339
			"000000000000000000000000000000000000",	-- 524 - 340
			"000000000000000000000000000000000000",	-- 525 - 341
			"000000000000000000000000000000000000",	-- 526 - 342
			"000000000000000000000000000000000000",	-- 527 - 343
			"000000000000000000000000000000000000",	-- 530 - 344
			"000000000000000000000000000000000000",	-- 531 - 345
			"000000000000000000000000000000000000",	-- 532 - 346
			"000000000000000000000000000000000000",	-- 533 - 347
			"000000000000000000000000000000000000",	-- 534 - 348
			"000000000000000000000000000000000000",	-- 535 - 349
			"000000000000000000000000000000000000",	-- 536 - 350
			"000000000000000000000000000000000000",	-- 537 - 351
			"000000000000000000000000000000000000",	-- 540 - 352
			"000000000000000000000000000000000000",	-- 541 - 353
			"000000000000000000000000000000000000",	-- 542 - 354
			"000000000000000000000000000000000000",	-- 543 - 355
			"000000000000000000000000000000000000",	-- 544 - 356
			"000000000000000000000000000000000000",	-- 545 - 357
			"000000000000000000000000000000000000",	-- 546 - 358
			"000000000000000000000000000000000000",	-- 547 - 359
			"000000000000000000000000000000000000",	-- 550 - 360
			"000000000000000000000000000000000000",	-- 551 - 361
			"000000000000000000000000000000000000",	-- 552 - 362
			"000000000000000000000000000000000000",	-- 553 - 363
			"000000000000000000000000000000000000",	-- 554 - 364
			"000000000000000000000000000000000000",	-- 555 - 365
			"000000000000000000000000000000000000",	-- 556 - 366
			"000000000000000000000000000000000000",	-- 557 - 367
			"000000000000000000000000000000000000",	-- 560 - 368
			"000000000000000000000000000000000000",	-- 561 - 369
			"000000000000000000000000000000000000",	-- 562 - 370
			"000000000000000000000000000000000000",	-- 563 - 371
			"000000000000000000000000000000000000",	-- 564 - 372
			"000000000000000000000000000000000000",	-- 565 - 373
			"000000000000000000000000000000000000",	-- 566 - 374
			"000000000000000000000000000000000000",	-- 567 - 375
			"000000000000000000000000000000000000",	-- 570 - 376
			"000000000000000000000000000000000000",	-- 571 - 377
			"000000000000000000000000000000000000",	-- 572 - 378
			"000000000000000000000000000000000000",	-- 573 - 379
			"000000000000000000000000000000000000",	-- 574 - 380
			"000000000000000000000000000000000000",	-- 575 - 381
			"000000000000000000000000000000000000",	-- 576 - 382
			"000000000000000000000000000000000000",	-- 577 - 383
			"110000001110100000000000000000110000",	-- 600 - 384
			"110000010000000000000111000000000000",	-- 601 - 385
			"110000011001111101000000000000000000",	-- 602 - 386
			"110000100000100010000000100000000000",	-- 603 - 387
			"000000000101100100000000000001000001",	-- 604 - 388
			"000000000000000000000000000000000000",	-- 605 - 389
			"000000000000000000000000000000000000",	-- 606 - 390
			"000000000000000000000000000000000000",	-- 607 - 391
			"110001001110100001000010011010000000",	-- 610 - 392
			"110001010001111100000000000001000000",	-- 611 - 393
			"000000000001000100000000000000000001",	-- 612 - 394
			"000000000000000000000000000000000000",	-- 613 - 395
			"000000000000000000000000000000000000",	-- 614 - 396
			"000000000000000000000000000000000000",	-- 615 - 397
			"000000000000000000000000000000000000",	-- 616 - 398
			"000000000000000000000000000000000000",	-- 617 - 399
			"000000000101100100000000000000010000",	-- 620 - 400
			"000000000000000000000000000000000000",	-- 621 - 401
			"000000000000000000000000000000000000",	-- 622 - 402
			"000000000000000000000000000000000000",	-- 623 - 403
			"000000000000000000000000000000000000",	-- 624 - 404
			"000000000000000000000000000000000000",	-- 625 - 405
			"000000000000000000000000000000000000",	-- 626 - 406
			"000000000000000000000000000000000000",	-- 627 - 407
			"110011001110100001000010011011000000",	-- 630 - 408
			"110011010001000100000000000000000000",	-- 631 - 409
			"110011011001100001000010010010000000",	-- 632 - 410
			"110011100001111100000000000001000000",	-- 633 - 411
			"000000000001011000000000000000100001",	-- 634 - 412
			"000000000000000000000000000000000000",	-- 635 - 413
			"000000000000000000000000000000000000",	-- 636 - 414
			"000000000000000000000000000000000000",	-- 637 - 415
			"000000000000000000000000000000000000",	-- 640 - 416
			"000000000000000000000000000000000000",	-- 641 - 417
			"000000000000000000000000000000000000",	-- 642 - 418
			"000000000000000000000000000000000000",	-- 643 - 419
			"000000000000000000000000000000000000",	-- 644 - 420
			"000000000000000000000000000000000000",	-- 645 - 421
			"000000000000000000000000000000000000",	-- 646 - 422
			"000000000000000000000000000000000000",	-- 647 - 423
			"000000000000000000000000000000000000",	-- 650 - 424
			"000000000000000000000000000000000000",	-- 651 - 425
			"000000000000000000000000000000000000",	-- 652 - 426
			"000000000000000000000000000000000000",	-- 653 - 427
			"000000000000000000000000000000000000",	-- 654 - 428
			"000000000000000000000000000000000000",	-- 655 - 429
			"000000000000000000000000000000000000",	-- 656 - 430
			"000000000000000000000000000000000000",	-- 657 - 431
			"000000000000000000000000000000000000",	-- 660 - 432
			"000000000000000000000000000000000000",	-- 661 - 433
			"000000000000000000000000000000000000",	-- 662 - 434
			"000000000000000000000000000000000000",	-- 663 - 435
			"000000000000000000000000000000000000",	-- 664 - 436
			"000000000000000000000000000000000000",	-- 665 - 437
			"000000000000000000000000000000000000",	-- 666 - 438
			"000000000000000000000000000000000000",	-- 667 - 439
			"000000000000000000000000000000000000",	-- 670 - 440
			"000000000000000000000000000000000000",	-- 671 - 441
			"000000000000000000000000000000000000",	-- 672 - 442
			"000000000000000000000000000000000000",	-- 673 - 443
			"000000000000000000000000000000000000",	-- 674 - 444
			"000000000000000000000000000000000000",	-- 675 - 445
			"000000000000000000000000000000000000",	-- 676 - 446
			"000000000000000000000000000000000000",	-- 677 - 447
			"111000001110100000000000000000110000",	-- 700 - 448
			"111000010000000000000111000000000000",	-- 701 - 449
			"111000011001100001000000000000110000",	-- 702 - 450
			"111000100110000010000111100001000000",	-- 703 - 451
			"111000101001111101000000000000000000",	-- 704 - 452
			"111000110000100010001111100001000000",	-- 705 - 453
			"000000000001100100000000000000000000",	-- 706 - 454
			"000000000000000000000000000000000000",	-- 707 - 455
			"000000000000000000000000000000000000",	-- 710 - 456
			"000000000000000000000000000000000000",	-- 711 - 457
			"000000000000000000000000000000000000",	-- 712 - 458
			"000000000000000000000000000000000000",	-- 713 - 459
			"000000000000000000000000000000000000",	-- 714 - 460
			"000000000000000000000000000000000000",	-- 715 - 461
			"000000000000000000000000000000000000",	-- 716 - 462
			"000000000000000000000000000000000000",	-- 717 - 463
			"000000000000000000000000000000000000",	-- 720 - 464
			"000000000000000000000000000000000000",	-- 721 - 465
			"000000000000000000000000000000000000",	-- 722 - 466
			"000000000000000000000000000000000000",	-- 723 - 467
			"000000000000000000000000000000000000",	-- 724 - 468
			"000000000000000000000000000000000000",	-- 725 - 469
			"000000000000000000000000000000000000",	-- 726 - 470
			"000000000000000000000000000000000000",	-- 727 - 471
			"000000000000000000000000000000000000",	-- 730 - 472
			"000000000000000000000000000000000000",	-- 731 - 473
			"000000000000000000000000000000000000",	-- 732 - 474
			"000000000000000000000000000000000000",	-- 733 - 475
			"000000000000000000000000000000000000",	-- 734 - 476
			"000000000000000000000000000000000000",	-- 735 - 477
			"000000000000000000000000000000000000",	-- 736 - 478
			"000000000000000000000000000000000000",	-- 737 - 479
			"000000000000000000000000000000000000",	-- 740 - 480
			"000000000000000000000000000000000000",	-- 741 - 481
			"000000000000000000000000000000000000",	-- 742 - 482
			"000000000000000000000000000000000000",	-- 743 - 483
			"000000000000000000000000000000000000",	-- 744 - 484
			"000000000000000000000000000000000000",	-- 745 - 485
			"000000000000000000000000000000000000",	-- 746 - 486
			"000000000000000000000000000000000000",	-- 747 - 487
			"000000000000000000000000000000000000",	-- 750 - 488
			"000000000000000000000000000000000000",	-- 751 - 489
			"000000000000000000000000000000000000",	-- 752 - 490
			"000000000000000000000000000000000000",	-- 753 - 491
			"000000000000000000000000000000000000",	-- 754 - 492
			"000000000000000000000000000000000000",	-- 755 - 493
			"000000000000000000000000000000000000",	-- 756 - 494
			"000000000000000000000000000000000000",	-- 757 - 495
			"000000000000000000000000000000000000",	-- 760 - 496
			"000000000000000000000000000000000000",	-- 761 - 497
			"000000000000000000000000000000000000",	-- 762 - 498
			"000000000000000000000000000000000000",	-- 763 - 499
			"000000000000000000000000000000000000",	-- 764 - 500
			"000000000000000000000000000000000000",	-- 765 - 501
			"000000000000000000000000000000000000",	-- 766 - 502
			"000000000000000000000000000000000000",	-- 767 - 503
			"000000000000000000000000000000000000",	-- 770 - 504
			"000000000000000000000000000000000000",	-- 771 - 505
			"000000000000000000000000000000000000",	-- 772 - 506
			"000000000000000000000000000000000000",	-- 773 - 507
			"000000000000000000000000000000000000",	-- 774 - 508
			"000000000000000000000000000000000000",	-- 775 - 509
			"000000000000000000000000000000000000",	-- 776 - 510
			"000000000000000000000000000000000000"	-- 777 - 511			
    );
begin
 
	process(clock) is
	begin
			if(start_signal = '1') then
					data_output <= mem(8#510#); -- At starting the processor make one NOP
			elsif(rising_edge(clock)) then
					data_output <= mem(conv_integer(unsigned(address)));
			end if;
	end process;
 
end a_code_store_rom;